library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_textio.all;

library std;
use std.textio.all;

entity data_maker is  
  port (
    CLK     : in  std_logic;
    RST_n   : in  std_logic;
    VOUT    : out std_logic;
    DOUT    : out std_logic_vector(12 downto 0);
    H0      : out std_logic_vector(12 downto 0); --coefficients
    H1      : out std_logic_vector(12 downto 0);
    H2      : out std_logic_vector(12 downto 0);
   -- H3      : out std_logic_vector(12 downto 0);
    END_SIM : out std_logic);
end data_maker;

architecture beh of data_maker is

  constant tco : time := 1 ns;
  --signal k: std_logic_vector(12 downto 0);
  signal sEndSim : std_logic;
  signal END_SIM_i : std_logic_vector(0 to 10); 
  signal svalid: std_logic; --user signal 
  signal sx: std_logic_vector(12 downto 0);
  signal SDOUT:std_logic_vector(12 downto 0);
  
begin  -- beh
 -- k<=conv_std_logic_vector(1265,13);
  H0 <= conv_std_logic_vector(-649,13); --a1
  H1 <= conv_std_logic_vector(1723,13); --b0
  H2 <= conv_std_logic_vector(1723,13); --b1
 -- H3 <= conv_std_logic_vector(9151,12);  

  process (CLK, RST_n)
    file fp_in : text open READ_MODE is "./matlab_VIN/samples.txt"; --change path
    variable line_in : line;
    variable k: integer:=666;
    --variable sx: integer;
    variable x : integer;
  begin  -- process
    if RST_n = '0' then                 -- asynchronous reset (active low)
      DOUT <= (others => '0') after tco;      
      VOUT <= '0' after tco;
      sEndSim <= '0' after tco;
    elsif CLK'event and CLK = '1' then  -- rising clock edge
      if not endfile(fp_in) then
        readline(fp_in, line_in);
        read(line_in, x);
		--sx<=conv_std_logic_vector(x, 13);
		if(x=k) then 
		VOUT <= '0' after tco;
      sEndSim <= '0' after tco;
      
		else
       	DOUT <= conv_std_logic_vector(x, 13) after tco;
        VOUT <= '1' after tco;
        sEndSim <= '0' after tco;
		end if;
      else
        VOUT <= '0' after tco;        
        sEndSim <= '1' after tco;
      end if;
    end if;
  end process;

  process (CLK, RST_n) --after 10 Vout=0 it stops the simulation
  begin  -- process
    if RST_n = '0' then                 -- asynchronous reset (active low)
      END_SIM_i <= (others => '0') after tco;
    elsif CLK'event and CLK = '1' then  -- rising clock edge
      END_SIM_i(0) <= sEndSim after tco;
      END_SIM_i(1 to 10) <= END_SIM_i(0 to 9) after tco;
    end if;
  end process;



          

  END_SIM <= END_SIM_i(10);  

end beh;
