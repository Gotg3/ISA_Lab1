library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


package filter_package is

	constant nb: integer:=13; --parallelism of the filter
	constant  N:  integer:=1;	 --order of the filter
	
end package filter_package;